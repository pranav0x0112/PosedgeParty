interface intf();
  logic d;
  logic clk;
  logic q;
  
endinterface	